parameter DIN_WIDTH = 18;
parameter COEFF_WIDTH = 16;
parameter DOUT_WIDTH = 31;
parameter NUM_CHN = 2;
parameter NUM_FACTOR = 1;
parameter TAPS_SIZE = 22;
parameter NUM_TDM = 1;
parameter COEFF_PATH = "./coeff.dat";
